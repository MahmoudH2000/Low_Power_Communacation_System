module moduleName #(
    parameter width = 8
) (
    // input & outputs ports
    
);
    
endmodule