module Rx_control (
    // input & output ports
    
);
    
endmodule